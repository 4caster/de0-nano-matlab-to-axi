
module pd_file (
	clk_clk,
	reset_reset_n,
	ledr_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	ledr_export;
endmodule

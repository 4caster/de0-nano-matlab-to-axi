-- pd_file.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pd_file is
	port (
		clk_clk       : in  std_logic                    := '0'; --   clk.clk
		ledr_export   : out std_logic_vector(7 downto 0);        --  ledr.export
		reset_reset_n : in  std_logic                    := '0'  -- reset.reset_n
	);
end entity pd_file;

architecture rtl of pd_file is
	component hdlverifier_axi_master is
		generic (
			JTAG_ID        : integer := 56;
			ID_WIDTH       : integer := 1;
			AXI_DATA_WIDTH : integer := 32;
			AXI_ADDR_WIDTH : integer := 32
		);
		port (
			axi4m_awaddr  : out std_logic_vector(31 downto 0);                    -- awaddr
			axi4m_awprot  : out std_logic_vector(2 downto 0);                     -- awprot
			axi4m_awvalid : out std_logic;                                        -- awvalid
			axi4m_awready : in  std_logic                     := 'X';             -- awready
			axi4m_wdata   : out std_logic_vector(31 downto 0);                    -- wdata
			axi4m_wlast   : out std_logic;                                        -- wlast
			axi4m_wvalid  : out std_logic;                                        -- wvalid
			axi4m_wready  : in  std_logic                     := 'X';             -- wready
			axi4m_bvalid  : in  std_logic                     := 'X';             -- bvalid
			axi4m_bready  : out std_logic;                                        -- bready
			axi4m_araddr  : out std_logic_vector(31 downto 0);                    -- araddr
			axi4m_arprot  : out std_logic_vector(2 downto 0);                     -- arprot
			axi4m_arvalid : out std_logic;                                        -- arvalid
			axi4m_arready : in  std_logic                     := 'X';             -- arready
			axi4m_rdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			axi4m_rvalid  : in  std_logic                     := 'X';             -- rvalid
			axi4m_rready  : out std_logic;                                        -- rready
			axi4m_arburst : out std_logic_vector(1 downto 0);                     -- arburst
			axi4m_arcache : out std_logic_vector(3 downto 0);                     -- arcache
			axi4m_arlen   : out std_logic_vector(7 downto 0);                     -- arlen
			axi4m_arlock  : out std_logic;                                        -- arlock
			axi4m_arqos   : out std_logic_vector(3 downto 0);                     -- arqos
			axi4m_arsize  : out std_logic_vector(2 downto 0);                     -- arsize
			axi4m_awburst : out std_logic_vector(1 downto 0);                     -- awburst
			axi4m_awcache : out std_logic_vector(3 downto 0);                     -- awcache
			axi4m_awid    : out std_logic_vector(0 downto 0);                     -- awid
			axi4m_awlen   : out std_logic_vector(7 downto 0);                     -- awlen
			axi4m_awlock  : out std_logic;                                        -- awlock
			axi4m_awqos   : out std_logic_vector(3 downto 0);                     -- awqos
			axi4m_awsize  : out std_logic_vector(2 downto 0);                     -- awsize
			axi4m_bresp   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			axi4m_rid     : in  std_logic                     := 'X';             -- rid
			axi4m_rlast   : in  std_logic                     := 'X';             -- rlast
			axi4m_rresp   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			axi4m_wstrb   : out std_logic_vector(3 downto 0);                     -- wstrb
			axi4m_arid    : out std_logic_vector(0 downto 0);                     -- arid
			axi4m_bid     : in  std_logic                     := 'X';             -- bid
			aclk          : in  std_logic                     := 'X';             -- clk
			aresetn       : in  std_logic                     := 'X'              -- reset_n
		);
	end component hdlverifier_axi_master;

	component pd_file_ledr is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component pd_file_ledr;

	component pd_file_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component pd_file_onchip_memory2_0;

	component pd_file_mm_interconnect_0 is
		port (
			MATLAB_as_AXI_Master_0_axm_m0_awid                         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- awid
			MATLAB_as_AXI_Master_0_axm_m0_awaddr                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			MATLAB_as_AXI_Master_0_axm_m0_awlen                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			MATLAB_as_AXI_Master_0_axm_m0_awsize                       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			MATLAB_as_AXI_Master_0_axm_m0_awburst                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			MATLAB_as_AXI_Master_0_axm_m0_awlock                       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- awlock
			MATLAB_as_AXI_Master_0_axm_m0_awcache                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			MATLAB_as_AXI_Master_0_axm_m0_awprot                       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			MATLAB_as_AXI_Master_0_axm_m0_awqos                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awqos
			MATLAB_as_AXI_Master_0_axm_m0_awvalid                      : in  std_logic                     := 'X';             -- awvalid
			MATLAB_as_AXI_Master_0_axm_m0_awready                      : out std_logic;                                        -- awready
			MATLAB_as_AXI_Master_0_axm_m0_wdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			MATLAB_as_AXI_Master_0_axm_m0_wstrb                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			MATLAB_as_AXI_Master_0_axm_m0_wlast                        : in  std_logic                     := 'X';             -- wlast
			MATLAB_as_AXI_Master_0_axm_m0_wvalid                       : in  std_logic                     := 'X';             -- wvalid
			MATLAB_as_AXI_Master_0_axm_m0_wready                       : out std_logic;                                        -- wready
			MATLAB_as_AXI_Master_0_axm_m0_bid                          : out std_logic_vector(0 downto 0);                     -- bid
			MATLAB_as_AXI_Master_0_axm_m0_bresp                        : out std_logic_vector(1 downto 0);                     -- bresp
			MATLAB_as_AXI_Master_0_axm_m0_bvalid                       : out std_logic;                                        -- bvalid
			MATLAB_as_AXI_Master_0_axm_m0_bready                       : in  std_logic                     := 'X';             -- bready
			MATLAB_as_AXI_Master_0_axm_m0_arid                         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- arid
			MATLAB_as_AXI_Master_0_axm_m0_araddr                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			MATLAB_as_AXI_Master_0_axm_m0_arlen                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			MATLAB_as_AXI_Master_0_axm_m0_arsize                       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			MATLAB_as_AXI_Master_0_axm_m0_arburst                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			MATLAB_as_AXI_Master_0_axm_m0_arlock                       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- arlock
			MATLAB_as_AXI_Master_0_axm_m0_arcache                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			MATLAB_as_AXI_Master_0_axm_m0_arprot                       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			MATLAB_as_AXI_Master_0_axm_m0_arqos                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arqos
			MATLAB_as_AXI_Master_0_axm_m0_arvalid                      : in  std_logic                     := 'X';             -- arvalid
			MATLAB_as_AXI_Master_0_axm_m0_arready                      : out std_logic;                                        -- arready
			MATLAB_as_AXI_Master_0_axm_m0_rid                          : out std_logic_vector(0 downto 0);                     -- rid
			MATLAB_as_AXI_Master_0_axm_m0_rdata                        : out std_logic_vector(31 downto 0);                    -- rdata
			MATLAB_as_AXI_Master_0_axm_m0_rresp                        : out std_logic_vector(1 downto 0);                     -- rresp
			MATLAB_as_AXI_Master_0_axm_m0_rlast                        : out std_logic;                                        -- rlast
			MATLAB_as_AXI_Master_0_axm_m0_rvalid                       : out std_logic;                                        -- rvalid
			MATLAB_as_AXI_Master_0_axm_m0_rready                       : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			MATLAB_as_AXI_Master_0_aresetn_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			ledr_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			ledr_s1_write                                              : out std_logic;                                        -- write
			ledr_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ledr_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			ledr_s1_chipselect                                         : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_address                                : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                  : out std_logic                                         -- clken
		);
	end component pd_file_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal matlab_as_axi_master_0_axm_m0_awburst            : std_logic_vector(1 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awburst -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awburst
	signal matlab_as_axi_master_0_axm_m0_arlen              : std_logic_vector(7 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arlen -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arlen
	signal matlab_as_axi_master_0_axm_m0_arqos              : std_logic_vector(3 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arqos -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arqos
	signal matlab_as_axi_master_0_axm_m0_wready             : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_wready -> MATLAB_as_AXI_Master_0:axi4m_wready
	signal matlab_as_axi_master_0_axm_m0_wstrb              : std_logic_vector(3 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_wstrb -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_wstrb
	signal matlab_as_axi_master_0_axm_m0_rid                : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rid -> MATLAB_as_AXI_Master_0:axi4m_rid
	signal matlab_as_axi_master_0_axm_m0_rready             : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_rready -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rready
	signal matlab_as_axi_master_0_axm_m0_awlen              : std_logic_vector(7 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awlen -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awlen
	signal matlab_as_axi_master_0_axm_m0_awqos              : std_logic_vector(3 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awqos -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awqos
	signal matlab_as_axi_master_0_axm_m0_arcache            : std_logic_vector(3 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arcache -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arcache
	signal matlab_as_axi_master_0_axm_m0_wvalid             : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_wvalid -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_wvalid
	signal matlab_as_axi_master_0_axm_m0_araddr             : std_logic_vector(31 downto 0); -- MATLAB_as_AXI_Master_0:axi4m_araddr -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_araddr
	signal matlab_as_axi_master_0_axm_m0_arprot             : std_logic_vector(2 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arprot -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arprot
	signal matlab_as_axi_master_0_axm_m0_awprot             : std_logic_vector(2 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awprot -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awprot
	signal matlab_as_axi_master_0_axm_m0_wdata              : std_logic_vector(31 downto 0); -- MATLAB_as_AXI_Master_0:axi4m_wdata -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_wdata
	signal matlab_as_axi_master_0_axm_m0_arvalid            : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_arvalid -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arvalid
	signal matlab_as_axi_master_0_axm_m0_awcache            : std_logic_vector(3 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awcache -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awcache
	signal matlab_as_axi_master_0_axm_m0_arid               : std_logic_vector(0 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arid -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arid
	signal matlab_as_axi_master_0_axm_m0_arlock             : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_arlock -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arlock
	signal matlab_as_axi_master_0_axm_m0_awlock             : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_awlock -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awlock
	signal matlab_as_axi_master_0_axm_m0_awaddr             : std_logic_vector(31 downto 0); -- MATLAB_as_AXI_Master_0:axi4m_awaddr -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awaddr
	signal matlab_as_axi_master_0_axm_m0_arready            : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arready -> MATLAB_as_AXI_Master_0:axi4m_arready
	signal matlab_as_axi_master_0_axm_m0_bresp              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_bresp -> MATLAB_as_AXI_Master_0:axi4m_bresp
	signal matlab_as_axi_master_0_axm_m0_rdata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rdata -> MATLAB_as_AXI_Master_0:axi4m_rdata
	signal matlab_as_axi_master_0_axm_m0_awready            : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awready -> MATLAB_as_AXI_Master_0:axi4m_awready
	signal matlab_as_axi_master_0_axm_m0_arburst            : std_logic_vector(1 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arburst -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arburst
	signal matlab_as_axi_master_0_axm_m0_arsize             : std_logic_vector(2 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_arsize -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_arsize
	signal matlab_as_axi_master_0_axm_m0_bready             : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_bready -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_bready
	signal matlab_as_axi_master_0_axm_m0_rlast              : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rlast -> MATLAB_as_AXI_Master_0:axi4m_rlast
	signal matlab_as_axi_master_0_axm_m0_wlast              : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_wlast -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_wlast
	signal matlab_as_axi_master_0_axm_m0_rresp              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rresp -> MATLAB_as_AXI_Master_0:axi4m_rresp
	signal matlab_as_axi_master_0_axm_m0_awid               : std_logic_vector(0 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awid -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awid
	signal matlab_as_axi_master_0_axm_m0_bid                : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_bid -> MATLAB_as_AXI_Master_0:axi4m_bid
	signal matlab_as_axi_master_0_axm_m0_bvalid             : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_bvalid -> MATLAB_as_AXI_Master_0:axi4m_bvalid
	signal matlab_as_axi_master_0_axm_m0_awvalid            : std_logic;                     -- MATLAB_as_AXI_Master_0:axi4m_awvalid -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awvalid
	signal matlab_as_axi_master_0_axm_m0_rvalid             : std_logic;                     -- mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_rvalid -> MATLAB_as_AXI_Master_0:axi4m_rvalid
	signal matlab_as_axi_master_0_axm_m0_awsize             : std_logic_vector(2 downto 0);  -- MATLAB_as_AXI_Master_0:axi4m_awsize -> mm_interconnect_0:MATLAB_as_AXI_Master_0_axm_m0_awsize
	signal mm_interconnect_0_ledr_s1_chipselect             : std_logic;                     -- mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	signal mm_interconnect_0_ledr_s1_readdata               : std_logic_vector(31 downto 0); -- ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	signal mm_interconnect_0_ledr_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ledr_s1_address -> ledr:address
	signal mm_interconnect_0_ledr_s1_write                  : std_logic;                     -- mm_interconnect_0:ledr_s1_write -> mm_interconnect_0_ledr_s1_write:in
	signal mm_interconnect_0_ledr_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata   : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address    : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write      : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken      : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal rst_controller_reset_out_reset                   : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:MATLAB_as_AXI_Master_0_aresetn_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req               : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                          : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_ledr_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_ledr_s1_write:inv -> ledr:write_n
	signal rst_controller_reset_out_reset_ports_inv         : std_logic;                     -- rst_controller_reset_out_reset:inv -> [MATLAB_as_AXI_Master_0:aresetn, ledr:reset_n]

begin

	matlab_as_axi_master_0 : component hdlverifier_axi_master
		generic map (
			JTAG_ID        => 56,
			ID_WIDTH       => 1,
			AXI_DATA_WIDTH => 32,
			AXI_ADDR_WIDTH => 32
		)
		port map (
			axi4m_awaddr  => matlab_as_axi_master_0_axm_m0_awaddr,     --  axm_m0.awaddr
			axi4m_awprot  => matlab_as_axi_master_0_axm_m0_awprot,     --        .awprot
			axi4m_awvalid => matlab_as_axi_master_0_axm_m0_awvalid,    --        .awvalid
			axi4m_awready => matlab_as_axi_master_0_axm_m0_awready,    --        .awready
			axi4m_wdata   => matlab_as_axi_master_0_axm_m0_wdata,      --        .wdata
			axi4m_wlast   => matlab_as_axi_master_0_axm_m0_wlast,      --        .wlast
			axi4m_wvalid  => matlab_as_axi_master_0_axm_m0_wvalid,     --        .wvalid
			axi4m_wready  => matlab_as_axi_master_0_axm_m0_wready,     --        .wready
			axi4m_bvalid  => matlab_as_axi_master_0_axm_m0_bvalid,     --        .bvalid
			axi4m_bready  => matlab_as_axi_master_0_axm_m0_bready,     --        .bready
			axi4m_araddr  => matlab_as_axi_master_0_axm_m0_araddr,     --        .araddr
			axi4m_arprot  => matlab_as_axi_master_0_axm_m0_arprot,     --        .arprot
			axi4m_arvalid => matlab_as_axi_master_0_axm_m0_arvalid,    --        .arvalid
			axi4m_arready => matlab_as_axi_master_0_axm_m0_arready,    --        .arready
			axi4m_rdata   => matlab_as_axi_master_0_axm_m0_rdata,      --        .rdata
			axi4m_rvalid  => matlab_as_axi_master_0_axm_m0_rvalid,     --        .rvalid
			axi4m_rready  => matlab_as_axi_master_0_axm_m0_rready,     --        .rready
			axi4m_arburst => matlab_as_axi_master_0_axm_m0_arburst,    --        .arburst
			axi4m_arcache => matlab_as_axi_master_0_axm_m0_arcache,    --        .arcache
			axi4m_arlen   => matlab_as_axi_master_0_axm_m0_arlen,      --        .arlen
			axi4m_arlock  => matlab_as_axi_master_0_axm_m0_arlock,     --        .arlock
			axi4m_arqos   => matlab_as_axi_master_0_axm_m0_arqos,      --        .arqos
			axi4m_arsize  => matlab_as_axi_master_0_axm_m0_arsize,     --        .arsize
			axi4m_awburst => matlab_as_axi_master_0_axm_m0_awburst,    --        .awburst
			axi4m_awcache => matlab_as_axi_master_0_axm_m0_awcache,    --        .awcache
			axi4m_awid    => matlab_as_axi_master_0_axm_m0_awid,       --        .awid
			axi4m_awlen   => matlab_as_axi_master_0_axm_m0_awlen,      --        .awlen
			axi4m_awlock  => matlab_as_axi_master_0_axm_m0_awlock,     --        .awlock
			axi4m_awqos   => matlab_as_axi_master_0_axm_m0_awqos,      --        .awqos
			axi4m_awsize  => matlab_as_axi_master_0_axm_m0_awsize,     --        .awsize
			axi4m_bresp   => matlab_as_axi_master_0_axm_m0_bresp,      --        .bresp
			axi4m_rid     => matlab_as_axi_master_0_axm_m0_rid,        --        .rid
			axi4m_rlast   => matlab_as_axi_master_0_axm_m0_rlast,      --        .rlast
			axi4m_rresp   => matlab_as_axi_master_0_axm_m0_rresp,      --        .rresp
			axi4m_wstrb   => matlab_as_axi_master_0_axm_m0_wstrb,      --        .wstrb
			axi4m_arid    => matlab_as_axi_master_0_axm_m0_arid,       --        .arid
			axi4m_bid     => matlab_as_axi_master_0_axm_m0_bid,        --        .bid
			aclk          => clk_clk,                                  --    aclk.clk
			aresetn       => rst_controller_reset_out_reset_ports_inv  -- aresetn.reset_n
		);

	ledr : component pd_file_ledr
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_ledr_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ledr_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ledr_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ledr_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ledr_s1_readdata,        --                    .readdata
			out_port   => ledr_export                                -- external_connection.export
		);

	onchip_memory2_0 : component pd_file_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	mm_interconnect_0 : component pd_file_mm_interconnect_0
		port map (
			MATLAB_as_AXI_Master_0_axm_m0_awid                         => matlab_as_axi_master_0_axm_m0_awid,               --                        MATLAB_as_AXI_Master_0_axm_m0.awid
			MATLAB_as_AXI_Master_0_axm_m0_awaddr                       => matlab_as_axi_master_0_axm_m0_awaddr,             --                                                     .awaddr
			MATLAB_as_AXI_Master_0_axm_m0_awlen                        => matlab_as_axi_master_0_axm_m0_awlen,              --                                                     .awlen
			MATLAB_as_AXI_Master_0_axm_m0_awsize                       => matlab_as_axi_master_0_axm_m0_awsize,             --                                                     .awsize
			MATLAB_as_AXI_Master_0_axm_m0_awburst                      => matlab_as_axi_master_0_axm_m0_awburst,            --                                                     .awburst
			MATLAB_as_AXI_Master_0_axm_m0_awlock(0)                    => matlab_as_axi_master_0_axm_m0_awlock,             --                                                     .awlock
			MATLAB_as_AXI_Master_0_axm_m0_awcache                      => matlab_as_axi_master_0_axm_m0_awcache,            --                                                     .awcache
			MATLAB_as_AXI_Master_0_axm_m0_awprot                       => matlab_as_axi_master_0_axm_m0_awprot,             --                                                     .awprot
			MATLAB_as_AXI_Master_0_axm_m0_awqos                        => matlab_as_axi_master_0_axm_m0_awqos,              --                                                     .awqos
			MATLAB_as_AXI_Master_0_axm_m0_awvalid                      => matlab_as_axi_master_0_axm_m0_awvalid,            --                                                     .awvalid
			MATLAB_as_AXI_Master_0_axm_m0_awready                      => matlab_as_axi_master_0_axm_m0_awready,            --                                                     .awready
			MATLAB_as_AXI_Master_0_axm_m0_wdata                        => matlab_as_axi_master_0_axm_m0_wdata,              --                                                     .wdata
			MATLAB_as_AXI_Master_0_axm_m0_wstrb                        => matlab_as_axi_master_0_axm_m0_wstrb,              --                                                     .wstrb
			MATLAB_as_AXI_Master_0_axm_m0_wlast                        => matlab_as_axi_master_0_axm_m0_wlast,              --                                                     .wlast
			MATLAB_as_AXI_Master_0_axm_m0_wvalid                       => matlab_as_axi_master_0_axm_m0_wvalid,             --                                                     .wvalid
			MATLAB_as_AXI_Master_0_axm_m0_wready                       => matlab_as_axi_master_0_axm_m0_wready,             --                                                     .wready
			MATLAB_as_AXI_Master_0_axm_m0_bid(0)                       => matlab_as_axi_master_0_axm_m0_bid,                --                                                     .bid
			MATLAB_as_AXI_Master_0_axm_m0_bresp                        => matlab_as_axi_master_0_axm_m0_bresp,              --                                                     .bresp
			MATLAB_as_AXI_Master_0_axm_m0_bvalid                       => matlab_as_axi_master_0_axm_m0_bvalid,             --                                                     .bvalid
			MATLAB_as_AXI_Master_0_axm_m0_bready                       => matlab_as_axi_master_0_axm_m0_bready,             --                                                     .bready
			MATLAB_as_AXI_Master_0_axm_m0_arid                         => matlab_as_axi_master_0_axm_m0_arid,               --                                                     .arid
			MATLAB_as_AXI_Master_0_axm_m0_araddr                       => matlab_as_axi_master_0_axm_m0_araddr,             --                                                     .araddr
			MATLAB_as_AXI_Master_0_axm_m0_arlen                        => matlab_as_axi_master_0_axm_m0_arlen,              --                                                     .arlen
			MATLAB_as_AXI_Master_0_axm_m0_arsize                       => matlab_as_axi_master_0_axm_m0_arsize,             --                                                     .arsize
			MATLAB_as_AXI_Master_0_axm_m0_arburst                      => matlab_as_axi_master_0_axm_m0_arburst,            --                                                     .arburst
			MATLAB_as_AXI_Master_0_axm_m0_arlock(0)                    => matlab_as_axi_master_0_axm_m0_arlock,             --                                                     .arlock
			MATLAB_as_AXI_Master_0_axm_m0_arcache                      => matlab_as_axi_master_0_axm_m0_arcache,            --                                                     .arcache
			MATLAB_as_AXI_Master_0_axm_m0_arprot                       => matlab_as_axi_master_0_axm_m0_arprot,             --                                                     .arprot
			MATLAB_as_AXI_Master_0_axm_m0_arqos                        => matlab_as_axi_master_0_axm_m0_arqos,              --                                                     .arqos
			MATLAB_as_AXI_Master_0_axm_m0_arvalid                      => matlab_as_axi_master_0_axm_m0_arvalid,            --                                                     .arvalid
			MATLAB_as_AXI_Master_0_axm_m0_arready                      => matlab_as_axi_master_0_axm_m0_arready,            --                                                     .arready
			MATLAB_as_AXI_Master_0_axm_m0_rid(0)                       => matlab_as_axi_master_0_axm_m0_rid,                --                                                     .rid
			MATLAB_as_AXI_Master_0_axm_m0_rdata                        => matlab_as_axi_master_0_axm_m0_rdata,              --                                                     .rdata
			MATLAB_as_AXI_Master_0_axm_m0_rresp                        => matlab_as_axi_master_0_axm_m0_rresp,              --                                                     .rresp
			MATLAB_as_AXI_Master_0_axm_m0_rlast                        => matlab_as_axi_master_0_axm_m0_rlast,              --                                                     .rlast
			MATLAB_as_AXI_Master_0_axm_m0_rvalid                       => matlab_as_axi_master_0_axm_m0_rvalid,             --                                                     .rvalid
			MATLAB_as_AXI_Master_0_axm_m0_rready                       => matlab_as_axi_master_0_axm_m0_rready,             --                                                     .rready
			clk_0_clk_clk                                              => clk_clk,                                          --                                            clk_0_clk.clk
			MATLAB_as_AXI_Master_0_aresetn_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                   -- MATLAB_as_AXI_Master_0_aresetn_reset_bridge_in_reset.reset
			ledr_s1_address                                            => mm_interconnect_0_ledr_s1_address,                --                                              ledr_s1.address
			ledr_s1_write                                              => mm_interconnect_0_ledr_s1_write,                  --                                                     .write
			ledr_s1_readdata                                           => mm_interconnect_0_ledr_s1_readdata,               --                                                     .readdata
			ledr_s1_writedata                                          => mm_interconnect_0_ledr_s1_writedata,              --                                                     .writedata
			ledr_s1_chipselect                                         => mm_interconnect_0_ledr_s1_chipselect,             --                                                     .chipselect
			onchip_memory2_0_s1_address                                => mm_interconnect_0_onchip_memory2_0_s1_address,    --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                  => mm_interconnect_0_onchip_memory2_0_s1_write,      --                                                     .write
			onchip_memory2_0_s1_readdata                               => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --                                                     .readdata
			onchip_memory2_0_s1_writedata                              => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --                                                     .writedata
			onchip_memory2_0_s1_byteenable                             => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                             => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --                                                     .chipselect
			onchip_memory2_0_s1_clken                                  => mm_interconnect_0_onchip_memory2_0_s1_clken       --                                                     .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_ledr_s1_write_ports_inv <= not mm_interconnect_0_ledr_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of pd_file
